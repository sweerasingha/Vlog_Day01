//Module Name: TwoInputAndGate

module TwoInputAndGate(
    input IN1, IN2,
    output OUT
);

assign OUT= IN1&IN2;

endmodule
