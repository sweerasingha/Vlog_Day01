module multiplexer_03(
    input [1:0] SEL,
    input [3:0] A,
    input [3:0] B,
    input [3:0] C,
    input [3:0] D,

    output reg [3:0] OUT
);
    always @ (SEL or A or B or C or D) begin
        case(SEL)
            2'b00: OUT <= A;
            2'b01: OUT <= B;
            2'b10: OUT <= C;
            2'b11: OUT <= D;
        endcase
    end
endmodule
